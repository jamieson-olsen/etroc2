-- ETROC2 readout testbench
-- jamieson olsen <jamieson@fnal.gov>

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.etroc2_package.all;

entity testbench is
end testbench;

architecture testbench_arch of testbench is

component etroc2 is
port(
    clock: in std_logic;
    reset: in std_logic;
	l1acc: in std_logic;
    d:     in  tdc_data_array_16_16_type;
    q:     out pixel_data_type
  );
end component;

signal clock: std_logic := '0';
signal reset: std_logic := '1';
signal l1acc: std_logic := '0';
signal d: tdc_data_array_16_16_type;

begin

clock <= not clock after 12.5ns; -- 40MHz BX

reset <= '1', '0' after 47ns;

main: process

-- some helper procedures

procedure clr_all is
begin
    InitLoopR: for R in 15 downto 0 loop
        InitLoopC: for C in 15 downto 0 loop
            d(R)(C).valid <= '0';
            d(R)(C).toa <= (others=>'0');
            d(R)(C).tot <= (others=>'0');
            d(R)(C).cal <= (others=>'0');
        end loop InitLoopC;
    end loop InitLoopR;
end procedure;

procedure set_pixel (constant row,col,toa,tot,cal: in integer) is
begin
    d(row)(col).valid <= '1';
    d(row)(col).tot   <= std_logic_vector(to_unsigned(tot,9));
    d(row)(col).toa   <= std_logic_vector(to_unsigned(toa,10));
    d(row)(col).cal   <= std_logic_vector(to_unsigned(cal,10));
end procedure;

procedure clr_pixel (constant row,col: in integer) is
begin
    d(row)(col).valid <= '0';
    d(row)(col).toa   <= (others=>'0');
    d(row)(col).tot   <= (others=>'0');
    d(row)(col).cal   <= (others=>'0');
end procedure;

begin 

-- do a few events by hand, gets tedious fast, will soon need to read events from file
-- when making fake TDC hits be sure TOT value is above threshold or else it will not
-- be written into the circular buffer!

clr_all;

wait for 1000ns;

-- first event

wait until falling_edge(clock);
set_pixel(4, 3, 122, 45, 98);
set_pixel(12, 4, 74, 15, 12);
set_pixel(9, 9, 41, 12, 49);
set_pixel(1, 14, 23, 92, 98);
wait until falling_edge(clock);
clr_all;
wait for 25ns * L1ACC_OFFSET;
l1acc <= '1';
wait until falling_edge(clock);
l1acc <= '0';

wait for 1000ns;  

-- a high occupancy event

wait until falling_edge(clock);
set_pixel(6, 11,  0, 21,  0);
set_pixel(15, 0,  0, 22,  0);
set_pixel(12, 15, 0, 23,  0);
set_pixel(15, 15, 0, 18,  0);
set_pixel(11, 0,  0, 43,  0);
set_pixel(1, 7, 0, 16, 0);
set_pixel(2, 7, 0, 78, 0);
set_pixel(3, 7, 0, 12, 0);
set_pixel(4, 7, 0, 32, 0);
set_pixel(5, 7, 0, 23, 0);
set_pixel(6, 7, 0, 75, 0);
set_pixel(7, 7, 0, 76, 0);
set_pixel(8, 7, 0, 77, 0);
set_pixel(9, 7, 0, 90, 0);
set_pixel(10, 7, 0, 13, 0);
set_pixel(11, 7, 0, 14, 0);
set_pixel(12, 7, 0, 15, 0);
set_pixel(13, 7, 0, 19, 0);
set_pixel(14, 7, 0, 19, 0);
set_pixel(15, 7, 0, 23, 0);
set_pixel(4, 8, 0, 21, 0);
set_pixel(12, 12, 0, 56, 0);
set_pixel(9, 3, 0, 11, 0);
set_pixel(12, 1, 0, 47, 0);
wait until falling_edge(clock);
clr_all;
wait for 25ns * L1ACC_OFFSET;
l1acc <= '1';
wait until falling_edge(clock);
l1acc <= '0';

wait for 1000ns;  

-- now try back to back to back L1accepts

wait until falling_edge(clock);
set_pixel(6, 1, 106, 107, 108);
set_pixel(6, 2, 109, 110, 111);
set_pixel(6, 3, 112, 113, 114);
set_pixel(6, 4, 115, 116, 117);
set_pixel(6, 5, 118, 118, 120);
set_pixel(9, 1, 121, 122, 123);

wait until falling_edge(clock);
clr_all;
set_pixel(8, 5, 206, 207, 208);
set_pixel(8, 6, 209, 210, 211);
set_pixel(8, 7, 212, 213, 214);
set_pixel(8, 8, 215, 216, 217);

wait until falling_edge(clock);
clr_all;
set_pixel(2,  12, 0, 61, 0);
set_pixel(3,  11, 0, 62, 0);
set_pixel(7,   5, 0, 63, 0);
set_pixel(14, 13, 0, 64, 0);
set_pixel(13, 13, 0, 65, 0);
set_pixel(2,   5, 0, 66, 0);
set_pixel(4,  11, 0, 67, 0);

wait until falling_edge(clock);
clr_all;
wait for 25ns * (L1ACC_OFFSET -2) ;
l1acc <= '1';
wait until falling_edge(clock);
wait until falling_edge(clock);
wait until falling_edge(clock);
l1acc <= '0';

wait;
end process main;


DUT: etroc2
port map( clock => clock, reset => reset, l1acc => l1acc, d => d );

end testbench_arch;
